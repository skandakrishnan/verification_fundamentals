// Code your design here
module add(
  input [3:0] a,b,
  output [4:0] sum
);
  
  assign sum = a+b;
endmodule

